/*
 * Description: Top level for AXI-Stream + APB based JPEG Encoder + ISP
 * 
 *
 * Authored by: Robert Metchev / Raumzeit Technologies (robert@raumzeit.co)
 *
 * CERN Open Hardware Licence Version 2 - Permissive
 *
 * Copyright (C) 2024 Robert Metchev
 */
`ifndef __AXIS_JPEG_ENCODER_VH__ 
`define __AXIS_JPEG_ENCODER_VH__

`endif // __AXIS_JPEG_ENCODER_VH__
